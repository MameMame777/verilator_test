class testclass;
  function new();
  endfunction
  task class_diplay;
    $display("This is a task called from class");
  endtask
endclass
