  export "DPI-C"    task enable_test_sv;
  export "DPI-C"    task check_count_sv;
  import "DPI-C" context function void enable_test();
  import "DPI-C" context function void check_count();